`define TEST_DATA_LENGTH 4096
`define TEST_DATA '{ \
  8'h9f,8'ha4,8'h2d,8'h91,8'h61,8'he4,8'h6a,8'h2a, \
  8'ha4,8'hf4,8'h2f,8'hc3,8'h23,8'he9,8'hed,8'h40, \
  8'h10,8'h0f,8'h81,8'h3b,8'hb7,8'h92,8'h7e,8'h63, \
  8'hc7,8'h9a,8'hd9,8'h75,8'ha1,8'h4f,8'h84,8'h81, \
  8'h46,8'hdc,8'h3d,8'h2c,8'ha8,8'hc7,8'h1a,8'ha1, \
  8'h32,8'h78,8'h52,8'h82,8'h47,8'hc7,8'h5a,8'h13, \
  8'he6,8'hb4,8'h5a,8'hd1,8'h25,8'h53,8'h74,8'ha8, \
  8'h3a,8'h04,8'hbb,8'hf6,8'h74,8'hda,8'hda,8'h62, \
  8'h21,8'hfc,8'h5d,8'he5,8'h2e,8'he5,8'h4e,8'hb7, \
  8'hdb,8'h78,8'hdb,8'h0f,8'ha2,8'h96,8'hc9,8'h82, \
  8'h57,8'h47,8'hb6,8'hf1,8'he3,8'hc9,8'h7d,8'h85, \
  8'hf2,8'h31,8'h41,8'hdb,8'hbf,8'hbc,8'ha6,8'h1c, \
  8'h35,8'h25,8'h39,8'hed,8'h0a,8'h15,8'hee,8'h83, \
  8'h04,8'h73,8'h6f,8'hf1,8'hc8,8'ha0,8'h76,8'h2f, \
  8'h72,8'h5e,8'h2a,8'he4,8'h41,8'h1a,8'hf8,8'h00, \
  8'hfd,8'h75,8'h54,8'h48,8'h5c,8'h32,8'he6,8'hf6, \
  8'hf3,8'h36,8'h2b,8'h92,8'h69,8'h65,8'h0d,8'h44, \
  8'hb1,8'h2b,8'h14,8'h33,8'ha9,8'h36,8'h8d,8'h1e, \
  8'h18,8'h70,8'h11,8'h33,8'h9b,8'h53,8'h87,8'h44, \
  8'ha3,8'he0,8'h6b,8'h57,8'h4e,8'hd5,8'h87,8'h62, \
  8'h80,8'h58,8'h6b,8'hba,8'hca,8'h5b,8'hec,8'hba, \
  8'ha7,8'h18,8'h6c,8'hc2,8'h69,8'h1f,8'h2f,8'h05, \
  8'hab,8'h4c,8'hff,8'h51,8'hed,8'hb0,8'h73,8'h39, \
  8'hc9,8'h4c,8'h52,8'h92,8'h02,8'h88,8'h1c,8'h28, \
  8'h98,8'h9d,8'hba,8'h9e,8'h01,8'h41,8'h59,8'he2, \
  8'h69,8'h47,8'h38,8'hf6,8'h96,8'hdc,8'h94,8'ha3, \
  8'h3f,8'h1c,8'h77,8'ha6,8'h44,8'h27,8'ha8,8'h52, \
  8'hc0,8'h66,8'h7b,8'h88,8'hde,8'h37,8'hdf,8'h26, \
  8'h2f,8'hec,8'h7f,8'h9b,8'hd1,8'h59,8'hea,8'hd9, \
  8'h19,8'haa,8'he6,8'he0,8'hbb,8'h82,8'h2f,8'h2d, \
  8'hd1,8'hc8,8'h2f,8'h83,8'h57,8'h03,8'h14,8'h32, \
  8'h66,8'h56,8'h1f,8'h38,8'h86,8'h7a,8'he6,8'ha8, \
  8'h21,8'ha5,8'h01,8'hc1,8'h51,8'h31,8'h42,8'h88, \
  8'h87,8'h85,8'hc1,8'h61,8'ha6,8'heb,8'h42,8'h14, \
  8'hb2,8'hc3,8'hfb,8'h4e,8'hd9,8'ha4,8'hf4,8'h7e, \
  8'h86,8'h5e,8'h3c,8'h21,8'h6b,8'h9c,8'h79,8'hda, \
  8'hf2,8'hb9,8'h0f,8'h62,8'h62,8'h4e,8'h75,8'h83, \
  8'h88,8'ha0,8'h4a,8'h71,8'h02,8'hfa,8'h97,8'h69, \
  8'hf5,8'h00,8'h3f,8'h41,8'h61,8'h09,8'hf5,8'h2a, \
  8'hb4,8'h55,8'h82,8'hf9,8'hb0,8'hc9,8'h09,8'h1a, \
  8'hd9,8'hb0,8'h9c,8'h6f,8'h5b,8'hb8,8'hd9,8'h5f, \
  8'ha5,8'h19,8'h94,8'h69,8'h1c,8'h65,8'h32,8'hc3, \
  8'h13,8'hb6,8'hba,8'hdb,8'h28,8'h1f,8'h2b,8'he4, \
  8'h76,8'hee,8'h96,8'h0d,8'h29,8'heb,8'hb3,8'hc1, \
  8'h51,8'hf3,8'h5c,8'h41,8'h7b,8'h56,8'hbf,8'h16, \
  8'h92,8'h28,8'h31,8'h18,8'hf4,8'h7f,8'hf7,8'hfd, \
  8'h8d,8'hc5,8'h68,8'h2d,8'hd3,8'h26,8'h08,8'h35, \
  8'h9d,8'h96,8'hc4,8'h32,8'hbd,8'h43,8'h28,8'hcc, \
  8'he3,8'h7c,8'he5,8'h5d,8'h56,8'he5,8'had,8'ha4, \
  8'h9b,8'h3d,8'h96,8'h0c,8'h15,8'h12,8'hfe,8'hff, \
  8'h97,8'hbe,8'h80,8'h6a,8'h18,8'h2b,8'he9,8'h1d, \
  8'h27,8'hb3,8'h25,8'h55,8'ha2,8'hcd,8'hee,8'hac, \
  8'he4,8'h14,8'h88,8'h16,8'hcc,8'h8a,8'ha2,8'h54, \
  8'h86,8'h8d,8'hf3,8'hc9,8'h49,8'h87,8'h18,8'h04, \
  8'h52,8'hbe,8'he8,8'h0c,8'hdb,8'h39,8'hba,8'hd0, \
  8'h67,8'hf3,8'h41,8'hc9,8'hb4,8'h70,8'h08,8'h6f, \
  8'h2b,8'h36,8'h6c,8'hb4,8'hc9,8'h42,8'h07,8'he2, \
  8'he1,8'hd5,8'hd1,8'h92,8'h6d,8'hf8,8'hbd,8'hb9, \
  8'hef,8'hd0,8'h54,8'h5b,8'h92,8'hd3,8'h48,8'hf5, \
  8'hf2,8'h2b,8'h1c,8'h32,8'h7b,8'haa,8'hcf,8'hc1, \
  8'ha7,8'h0d,8'hb5,8'h30,8'h5d,8'hac,8'h10,8'h73, \
  8'h20,8'h15,8'h8e,8'hea,8'hd1,8'he7,8'hc6,8'h2e, \
  8'h2e,8'h1c,8'h79,8'hf0,8'h89,8'ha4,8'h9f,8'hbc, \
  8'h8c,8'hdd,8'h12,8'h57,8'hec,8'h8e,8'hbc,8'h25, \
  8'h80,8'hcf,8'hf9,8'h86,8'he2,8'h29,8'h03,8'ha1, \
  8'hcb,8'h1c,8'hb3,8'h5d,8'h3e,8'h58,8'h40,8'h6a, \
  8'h4a,8'h37,8'h8e,8'h17,8'hdb,8'h08,8'h2e,8'ha9, \
  8'h07,8'h41,8'h70,8'hdd,8'hae,8'h02,8'he4,8'he3, \
  8'h26,8'hc8,8'hbf,8'hae,8'h3f,8'hdd,8'h09,8'ha4, \
  8'h95,8'ha4,8'hc4,8'h8c,8'hb8,8'h1d,8'hfc,8'h05, \
  8'h4f,8'ha7,8'h85,8'h3a,8'hfd,8'h81,8'h00,8'h77, \
  8'h38,8'h77,8'h88,8'h7d,8'h9f,8'h46,8'h39,8'h9d, \
  8'hf3,8'h5f,8'h24,8'hd7,8'h4b,8'hc1,8'hbc,8'he9, \
  8'h3a,8'h1e,8'h6f,8'hcd,8'haf,8'he9,8'h85,8'hd0, \
  8'h73,8'h11,8'h90,8'h80,8'hb4,8'h91,8'h3a,8'h34, \
  8'h1c,8'h90,8'h5d,8'h3f,8'h5e,8'h7c,8'hbc,8'hde, \
  8'h57,8'h43,8'hba,8'h50,8'h90,8'h6f,8'h7c,8'ha1, \
  8'hb2,8'ha5,8'hb1,8'hd3,8'he9,8'h73,8'h64,8'h9e, \
  8'ha9,8'hb4,8'hd2,8'h12,8'h9d,8'h7d,8'h91,8'hfa, \
  8'h89,8'h9b,8'h50,8'h51,8'h7f,8'h68,8'h71,8'hb2, \
  8'h16,8'h80,8'h91,8'h0b,8'h71,8'h95,8'h21,8'h86, \
  8'hb0,8'h0a,8'h9f,8'he4,8'h49,8'h4a,8'hc9,8'h4f, \
  8'h12,8'hb2,8'h0d,8'h9b,8'h3c,8'h91,8'h91,8'hda, \
  8'he0,8'h35,8'h9f,8'h2b,8'hb3,8'hdd,8'h71,8'h74, \
  8'h65,8'h42,8'ha7,8'hf9,8'h6e,8'h5c,8'h6c,8'he0, \
  8'h38,8'hd0,8'h3e,8'hc0,8'h56,8'h0f,8'h06,8'h31, \
  8'h44,8'h17,8'h31,8'h4e,8'hcb,8'hc9,8'hc6,8'h2f, \
  8'h48,8'ha7,8'h34,8'h29,8'h63,8'hd7,8'ha7,8'h06, \
  8'h17,8'hf0,8'h14,8'he5,8'h9b,8'hcf,8'h0a,8'ha6, \
  8'h39,8'hac,8'h96,8'hea,8'ha1,8'hc9,8'h03,8'h28, \
  8'ha5,8'hd3,8'h5e,8'h0e,8'h21,8'h50,8'hc8,8'h1a, \
  8'h71,8'h53,8'he2,8'hbb,8'hd7,8'hc5,8'ha0,8'hf0, \
  8'hc4,8'h65,8'h93,8'h7d,8'h58,8'hb0,8'h56,8'h4f, \
  8'h37,8'hea,8'hc5,8'hec,8'hfb,8'hd5,8'h0a,8'hb2, \
  8'h00,8'h09,8'hdf,8'ha5,8'h25,8'hb0,8'h87,8'hb0, \
  8'h2f,8'h51,8'h9e,8'h43,8'he8,8'h34,8'h43,8'h78, \
  8'hf8,8'h4c,8'he5,8'h58,8'h41,8'h74,8'h5d,8'hcd, \
  8'h79,8'h5c,8'h4e,8'h27,8'h72,8'h3d,8'had,8'h22, \
  8'h1b,8'h04,8'hb1,8'h88,8'hc5,8'h37,8'h53,8'hc7, \
  8'ha7,8'hef,8'hc2,8'h76,8'hbc,8'h08,8'h6d,8'hb5, \
  8'h4b,8'h58,8'hb0,8'hfe,8'h66,8'h72,8'h4a,8'hd1, \
  8'hca,8'ha8,8'h4f,8'hb1,8'h8c,8'ha5,8'h56,8'h6e, \
  8'hb1,8'h96,8'h68,8'hba,8'h66,8'h4f,8'h4c,8'h83, \
  8'hef,8'h0d,8'hce,8'h79,8'hb4,8'h15,8'h73,8'hd7, \
  8'h46,8'hd3,8'hc8,8'hc2,8'heb,8'h7a,8'h1e,8'h60, \
  8'h6b,8'h49,8'h1a,8'h0a,8'hbf,8'he0,8'ha8,8'h34, \
  8'h33,8'ha0,8'h38,8'h26,8'h68,8'h6c,8'h8e,8'h37, \
  8'hf0,8'h0e,8'h42,8'hc1,8'hff,8'he6,8'h77,8'hd3, \
  8'h31,8'hff,8'h6f,8'h3e,8'hb4,8'h0c,8'h2f,8'hba, \
  8'h7e,8'h0e,8'hf2,8'h61,8'hfa,8'h8b,8'h54,8'h82, \
  8'h0c,8'h32,8'h9d,8'h9c,8'h32,8'h12,8'h87,8'h8b, \
  8'h33,8'hfb,8'ha3,8'he5,8'h18,8'h98,8'h00,8'h20, \
  8'h25,8'h34,8'hf4,8'hbb,8'h8b,8'hfc,8'h93,8'hc5, \
  8'h02,8'h85,8'ha1,8'h03,8'h9b,8'h5a,8'h75,8'h93, \
  8'h76,8'h0e,8'h94,8'h58,8'hb7,8'h98,8'hdc,8'hb3, \
  8'h93,8'hb6,8'h87,8'h15,8'hc1,8'hfa,8'hec,8'h0b, \
  8'h06,8'h89,8'h42,8'h16,8'h04,8'hc2,8'h87,8'h86, \
  8'ha1,8'h7d,8'h47,8'hbb,8'h4f,8'hea,8'hbf,8'hfc, \
  8'h48,8'hc0,8'hc7,8'h50,8'hfa,8'ha6,8'hbf,8'hd2, \
  8'h5b,8'ha9,8'hd3,8'hc5,8'ha6,8'h02,8'h63,8'he7, \
  8'h17,8'h5b,8'h83,8'h00,8'h84,8'h98,8'haf,8'h9b, \
  8'ha1,8'h6b,8'h5a,8'hcb,8'hc4,8'h8e,8'hee,8'ha6, \
  8'hd9,8'hf6,8'h0c,8'h53,8'h33,8'h96,8'h5e,8'h35, \
  8'h0d,8'hba,8'h3e,8'h30,8'hc9,8'h8b,8'h4d,8'h6d, \
  8'h81,8'h21,8'hc5,8'hf4,8'hbd,8'h74,8'h53,8'hb3, \
  8'h41,8'h2b,8'h25,8'h87,8'h29,8'h65,8'h68,8'hc1, \
  8'hc3,8'hdb,8'hd1,8'hd8,8'h42,8'h3f,8'h79,8'hd5, \
  8'h5b,8'h87,8'h27,8'hca,8'h9c,8'hc8,8'hb8,8'hee, \
  8'h2f,8'hc5,8'h22,8'hdf,8'h50,8'heb,8'hed,8'h6e, \
  8'h0a,8'hae,8'hf1,8'h0c,8'hcd,8'h81,8'hf9,8'hd8, \
  8'h9e,8'h01,8'h79,8'hab,8'he2,8'h3c,8'h40,8'ha7, \
  8'hbf,8'h13,8'hcf,8'h91,8'h80,8'h65,8'h52,8'h63, \
  8'h42,8'h70,8'hbc,8'h3f,8'h70,8'h8e,8'hb9,8'h57, \
  8'hfb,8'h10,8'hf0,8'hfd,8'h8e,8'h5a,8'h12,8'h27, \
  8'h4d,8'h3c,8'h6a,8'ha2,8'hd3,8'hc2,8'hf0,8'hc0, \
  8'h7b,8'ha0,8'hfd,8'h80,8'h9e,8'hfb,8'hf2,8'hff, \
  8'h49,8'hda,8'h24,8'hd0,8'hce,8'hb2,8'he3,8'h8d, \
  8'hdf,8'hcb,8'h08,8'h31,8'hf6,8'hf4,8'hcc,8'h84, \
  8'h1d,8'h76,8'h37,8'ha1,8'hcd,8'h68,8'h3a,8'h02, \
  8'h01,8'he5,8'hb3,8'h4d,8'h8e,8'he2,8'hc7,8'h07, \
  8'h0d,8'h27,8'hf3,8'h2b,8'hd7,8'h32,8'h28,8'h51, \
  8'h8b,8'h9b,8'hc1,8'hf1,8'h4d,8'ha7,8'h20,8'h67, \
  8'h8c,8'h73,8'h1c,8'hc2,8'h3d,8'hf1,8'h90,8'h85, \
  8'hb4,8'h7d,8'h16,8'he7,8'h50,8'h9d,8'hb3,8'h40, \
  8'hef,8'h5f,8'h60,8'hcf,8'h5d,8'hbf,8'h46,8'h6d, \
  8'hb2,8'h45,8'hee,8'h8e,8'hef,8'hc3,8'h47,8'h44, \
  8'h2a,8'h8b,8'h10,8'h1e,8'ha3,8'h70,8'h89,8'heb, \
  8'h60,8'he9,8'hdc,8'hfd,8'h30,8'hc6,8'h92,8'h67, \
  8'hc0,8'h9a,8'hc7,8'h8a,8'h82,8'hff,8'h0c,8'hf5, \
  8'h79,8'h5f,8'h88,8'hbb,8'h4a,8'h21,8'hde,8'he0, \
  8'hdb,8'h2b,8'hb7,8'h07,8'hf2,8'hdc,8'h0a,8'h39, \
  8'h8d,8'hba,8'h90,8'h1a,8'h0a,8'ha1,8'h0d,8'hab, \
  8'h43,8'h29,8'h80,8'h4a,8'h02,8'h75,8'h72,8'h66, \
  8'h1d,8'he9,8'h81,8'h5f,8'ha2,8'h45,8'h1d,8'heb, \
  8'h05,8'h33,8'h5f,8'hb4,8'hf2,8'h35,8'hef,8'h8a, \
  8'h00,8'hdf,8'h84,8'h00,8'hee,8'hca,8'h10,8'he6, \
  8'ha8,8'h80,8'h9b,8'h0c,8'h56,8'he4,8'h9f,8'he5, \
  8'h13,8'he6,8'h49,8'hb5,8'hec,8'h7e,8'h76,8'h4c, \
  8'ha5,8'h31,8'hbd,8'h1b,8'h98,8'h72,8'h3a,8'h06, \
  8'hf0,8'h94,8'h39,8'hea,8'h2d,8'he0,8'h56,8'h6b, \
  8'h39,8'ha2,8'hdd,8'h9b,8'h5f,8'h4c,8'h06,8'h45, \
  8'h60,8'h85,8'h26,8'h5f,8'hdf,8'h47,8'h80,8'h7d, \
  8'he2,8'h30,8'ha4,8'h52,8'h7a,8'hc3,8'hc6,8'h59, \
  8'hf4,8'h54,8'he4,8'h0a,8'h6e,8'ha6,8'hec,8'hcb, \
  8'hee,8'hf6,8'hc2,8'hea,8'he1,8'hf1,8'h1e,8'h42, \
  8'h22,8'h5b,8'ha0,8'h86,8'h26,8'hc8,8'h46,8'hbd, \
  8'h14,8'h2c,8'hae,8'h56,8'h83,8'h0a,8'h75,8'h26, \
  8'hb3,8'h93,8'h09,8'h10,8'h87,8'hde,8'h19,8'hb5, \
  8'hdc,8'hf0,8'h04,8'h0b,8'h9a,8'h9f,8'hb0,8'hda, \
  8'h54,8'hc0,8'h0f,8'h28,8'h53,8'hbb,8'h01,8'h43, \
  8'h31,8'h6b,8'hda,8'hb6,8'hb6,8'h7e,8'hda,8'h34, \
  8'h62,8'hdc,8'h0a,8'h24,8'h1e,8'hd6,8'hc7,8'hdf, \
  8'he5,8'h78,8'h34,8'hc8,8'h42,8'h5f,8'h30,8'hdf, \
  8'h45,8'hc1,8'hbf,8'he6,8'h9d,8'h3e,8'h7d,8'h3f, \
  8'hea,8'h49,8'h0e,8'h0b,8'h49,8'hbe,8'h8f,8'hac, \
  8'h66,8'h86,8'h70,8'h27,8'he3,8'hb9,8'h64,8'h62, \
  8'hec,8'hf1,8'h73,8'hf2,8'hfe,8'h44,8'he3,8'h7d, \
  8'h83,8'h33,8'ha0,8'h9f,8'hbd,8'h67,8'h82,8'hf0, \
  8'h17,8'h4d,8'h61,8'h3a,8'h40,8'hc1,8'h24,8'hb7, \
  8'hf1,8'h3b,8'hd4,8'hc9,8'h9e,8'hfb,8'hd1,8'h96, \
  8'h9c,8'h28,8'hc2,8'hc3,8'h4b,8'h71,8'h00,8'h87, \
  8'hcc,8'h84,8'hda,8'h2e,8'hb4,8'hb5,8'h8b,8'hd0, \
  8'hc2,8'h85,8'h4d,8'h6c,8'hfb,8'h26,8'h92,8'ha3, \
  8'h2e,8'hb6,8'h6d,8'hb6,8'h72,8'hef,8'h85,8'h90, \
  8'h19,8'hbf,8'h39,8'hd9,8'h2e,8'hc0,8'hbb,8'h14, \
  8'hb6,8'h55,8'hf6,8'h8c,8'hcf,8'h9b,8'h2a,8'ha3, \
  8'hbb,8'h40,8'ha9,8'hb3,8'hda,8'h96,8'h15,8'h93, \
  8'h00,8'h63,8'h68,8'h64,8'h21,8'h83,8'hf0,8'h5b, \
  8'h88,8'h21,8'hba,8'h9c,8'h94,8'h97,8'h97,8'h04, \
  8'hbd,8'h81,8'h47,8'h60,8'hd1,8'h5c,8'h5a,8'h8d, \
  8'h4c,8'h9f,8'hfd,8'h52,8'h4d,8'he4,8'h28,8'h44, \
  8'h37,8'h3d,8'h76,8'hbb,8'h6f,8'hdc,8'h93,8'hf7, \
  8'h0c,8'h5d,8'h01,8'h4b,8'hc0,8'h5a,8'hea,8'hea, \
  8'h28,8'hc2,8'hca,8'h48,8'hd4,8'h4a,8'h19,8'h68, \
  8'h2b,8'h3b,8'hc0,8'h5a,8'h7a,8'hc9,8'h9a,8'h72, \
  8'hc6,8'hc6,8'hb8,8'h45,8'h76,8'h28,8'h67,8'he2, \
  8'h35,8'hbe,8'h3f,8'h95,8'h7f,8'h10,8'h11,8'h5b, \
  8'h40,8'h6c,8'he1,8'hc9,8'h0b,8'h92,8'h00,8'h02, \
  8'h41,8'hf7,8'hcb,8'h1f,8'h27,8'h48,8'hd2,8'h90, \
  8'h82,8'h50,8'h4e,8'hdc,8'h02,8'hf0,8'h35,8'hae, \
  8'h9f,8'h1e,8'h96,8'hfc,8'hab,8'hc5,8'h1a,8'h82, \
  8'h1b,8'h04,8'hb5,8'h36,8'h6b,8'h98,8'hc9,8'h4e, \
  8'h42,8'h8a,8'h9b,8'h3e,8'h11,8'h75,8'h11,8'haf, \
  8'he3,8'hc9,8'h2a,8'h0f,8'h36,8'h8e,8'hcc,8'h70, \
  8'h46,8'hdd,8'hde,8'h22,8'h3f,8'hf5,8'hc2,8'h98, \
  8'hee,8'h64,8'hd6,8'ha6,8'h46,8'h5d,8'hca,8'h6e, \
  8'ha0,8'h0c,8'he0,8'h43,8'hdb,8'h38,8'h50,8'ha4, \
  8'heb,8'he8,8'h06,8'he9,8'h2e,8'ha8,8'h78,8'h74, \
  8'hf6,8'h27,8'h68,8'hdc,8'h25,8'hb6,8'h49,8'h6a, \
  8'h0d,8'hf3,8'hf6,8'h61,8'h77,8'hda,8'h79,8'hcc, \
  8'hea,8'h8f,8'h74,8'hfc,8'h0e,8'h60,8'h50,8'hf9, \
  8'h26,8'h7b,8'h96,8'h28,8'hba,8'h9f,8'h82,8'h01, \
  8'h8e,8'he0,8'hca,8'h0e,8'hab,8'hbf,8'h19,8'h27, \
  8'hff,8'hd4,8'h86,8'h87,8'h1d,8'he4,8'hbe,8'h23, \
  8'h50,8'h60,8'hbb,8'hb8,8'hf5,8'h8e,8'h06,8'ha5, \
  8'h02,8'h18,8'h30,8'h5f,8'h58,8'hc5,8'h86,8'h09, \
  8'h8e,8'hd9,8'h47,8'h9d,8'h39,8'h25,8'hdb,8'h17, \
  8'h81,8'h71,8'h3e,8'hdc,8'h3b,8'ha3,8'h49,8'hc7, \
  8'h1d,8'h24,8'h79,8'h57,8'h72,8'he3,8'hcf,8'hfe, \
  8'hdd,8'h3a,8'h78,8'h3b,8'hac,8'hd9,8'h5a,8'hfd, \
  8'hb3,8'h7f,8'h6a,8'hda,8'h60,8'hd2,8'h84,8'h88, \
  8'hea,8'h34,8'h19,8'ha2,8'hea,8'hb8,8'hd3,8'h7e, \
  8'hc5,8'h24,8'h52,8'h35,8'h19,8'h7a,8'hcc,8'h13, \
  8'h85,8'h99,8'h09,8'h36,8'h60,8'hf0,8'h45,8'hb1, \
  8'hff,8'h45,8'he0,8'h08,8'h3c,8'hbc,8'hc2,8'h7b, \
  8'h28,8'h8a,8'hd4,8'h4c,8'h6d,8'h7e,8'hfe,8'hc1, \
  8'h68,8'h24,8'h7f,8'h13,8'ha2,8'hcf,8'hc8,8'h5e, \
  8'hd2,8'h03,8'h06,8'he3,8'hbd,8'h7a,8'hd1,8'h31, \
  8'hd8,8'hdb,8'h7c,8'ha6,8'h3e,8'h76,8'h83,8'h57, \
  8'h1a,8'h44,8'h6d,8'h37,8'h3c,8'heb,8'h19,8'h78, \
  8'h15,8'hbf,8'h57,8'hc3,8'hbe,8'h49,8'h96,8'h27, \
  8'h3a,8'hdc,8'h5c,8'hd7,8'h79,8'h92,8'hce,8'h8b, \
  8'h28,8'hb4,8'h8a,8'h58,8'h08,8'h06,8'ha1,8'h3d, \
  8'hb7,8'h73,8'h12,8'h01,8'h4c,8'h66,8'h9e,8'hdf, \
  8'hed,8'ha6,8'h2f,8'ha2,8'hbf,8'h5f,8'h26,8'h73, \
  8'hd3,8'h77,8'h54,8'hd0,8'hde,8'hb8,8'he2,8'hba, \
  8'h8b,8'h24,8'had,8'h04,8'hc9,8'h99,8'hbd,8'hf8, \
  8'h0a,8'hf5,8'h91,8'h72,8'ha3,8'h37,8'he5,8'h37, \
  8'h70,8'he8,8'hbf,8'h0f,8'h16,8'hac,8'h85,8'hd7, \
  8'hc1,8'h4f,8'h2a,8'h05,8'h7b,8'h94,8'hdd,8'hd4, \
  8'hf0,8'h5b,8'h51,8'h2a,8'h3b,8'h9a,8'hd2,8'h0a, \
  8'hb5,8'h39,8'hbd,8'hcc,8'ha1,8'h01,8'hb5,8'h8f, \
  8'hde,8'h18,8'h96,8'h00,8'h9b,8'h3f,8'h03,8'h51, \
  8'hf1,8'h3f,8'h3c,8'h35,8'h20,8'h05,8'h5b,8'h37, \
  8'hd2,8'hd1,8'h6e,8'h51,8'hfb,8'h2d,8'hbf,8'h7e, \
  8'h0d,8'h40,8'h14,8'ha7,8'h7c,8'h7f,8'hb8,8'h49, \
  8'hc2,8'h5e,8'h20,8'hd6,8'h20,8'h7f,8'hfe,8'h3d, \
  8'h09,8'hd5,8'h7a,8'hb8,8'h5e,8'h28,8'h58,8'ha0, \
  8'h90,8'hc9,8'he7,8'h93,8'h69,8'h3c,8'h7a,8'h75, \
  8'h58,8'h39,8'h32,8'h8f,8'h68,8'h46,8'hda,8'he0, \
  8'h70,8'hb9,8'h97,8'h4c,8'hea,8'h6b,8'h63,8'h97, \
  8'hbe,8'had,8'h2f,8'h44,8'h47,8'hd6,8'h9c,8'h84, \
  8'h62,8'hb2,8'h22,8'hc2,8'h98,8'h66,8'h63,8'h68, \
  8'hec,8'h50,8'hf9,8'hb5,8'h90,8'h54,8'ha8,8'hed, \
  8'h20,8'h23,8'h04,8'h5e,8'hcf,8'h60,8'h67,8'ha6, \
  8'h67,8'h59,8'hf6,8'h2e,8'he8,8'h01,8'ha3,8'h82, \
  8'h5c,8'h72,8'hac,8'h8c,8'h74,8'h39,8'h12,8'h96, \
  8'h1a,8'he8,8'h26,8'h59,8'h8f,8'hb6,8'h39,8'h79, \
  8'h2c,8'hff,8'hc1,8'hb8,8'he8,8'h62,8'h0a,8'hc8, \
  8'hdb,8'h72,8'hf1,8'hc7,8'h90,8'hfc,8'h90,8'h94, \
  8'h48,8'h96,8'h8f,8'he6,8'h3b,8'ha1,8'hfb,8'hd0, \
  8'h26,8'h2c,8'h34,8'hd2,8'h1d,8'h41,8'ha4,8'h1e, \
  8'h59,8'h63,8'hcd,8'h45,8'hd2,8'h32,8'h6b,8'hda, \
  8'hcb,8'h92,8'hbc,8'h93,8'h81,8'hd1,8'hd6,8'h08, \
  8'h14,8'hab,8'he3,8'h77,8'he5,8'h25,8'h8a,8'h5f, \
  8'h43,8'hc3,8'h02,8'h84,8'h85,8'h65,8'hc8,8'h08, \
  8'h81,8'he7,8'h4d,8'hc6,8'hc1,8'h92,8'h17,8'h80, \
  8'h34,8'hda,8'h88,8'hc4,8'hff,8'he3,8'hee,8'hd1, \
  8'h2f,8'hd0,8'h61,8'h63,8'hdb,8'h23,8'hc6,8'h55, \
  8'h41,8'he7,8'h90,8'h81,8'h7b,8'ha1,8'h62,8'h06, \
  8'h9b,8'h25,8'h2e,8'hf1,8'h1b,8'h0a,8'h2e,8'h95, \
  8'hff,8'hfd,8'h1a,8'h45,8'hb8,8'h78,8'h76,8'he2, \
  8'hdd,8'ha5,8'he9,8'hc6,8'h18,8'h60,8'ha5,8'h5e, \
  8'hd7,8'hdc,8'h99,8'h68,8'h0e,8'hd3,8'hb0,8'h42, \
  8'hc0,8'h8a,8'hff,8'h2a,8'h44,8'hf0,8'ha8,8'h8a, \
  8'h7a,8'hbd,8'h02,8'h9b,8'hfe,8'h01,8'hb9,8'h3c, \
  8'h65,8'h86,8'h12,8'h2a,8'h16,8'hdd,8'h11,8'h25, \
  8'h59,8'h65,8'h23,8'h89,8'hc8,8'hc2,8'ha8,8'h29, \
  8'he7,8'h48,8'h16,8'hf3,8'h94,8'h19,8'h3b,8'h13, \
  8'hda,8'hfc,8'h29,8'h6d,8'h44,8'h8d,8'h03,8'h98, \
  8'he2,8'h6c,8'h2b,8'hee,8'he3,8'h8c,8'hf2,8'h33, \
  8'h84,8'h07,8'h92,8'h65,8'h53,8'h7c,8'he8,8'h84, \
  8'h3f,8'h86,8'h7b,8'hda,8'h97,8'h34,8'hcd,8'h7f, \
  8'h2f,8'h22,8'hff,8'h7f,8'h25,8'ha3,8'h83,8'he7, \
  8'h2b,8'he5,8'h69,8'h1e,8'h4f,8'ha3,8'h32,8'h53, \
  8'he5,8'hb6,8'h33,8'ha5,8'hb4,8'he9,8'h70,8'hce, \
  8'hc0,8'hde,8'h93,8'hfa,8'h91,8'he5,8'ha0,8'hcf, \
  8'h7e,8'h80,8'hba,8'hc7,8'h1d,8'hb6,8'h0c,8'h5d, \
  8'h33,8'hc3,8'h98,8'h26,8'h68,8'hd4,8'h7c,8'hdb, \
  8'had,8'h33,8'he7,8'he8,8'h57,8'h97,8'hbf,8'hbc, \
  8'hcd,8'h31,8'h6e,8'hca,8'he3,8'h39,8'h8f,8'hff, \
  8'h12,8'h1d,8'hcf,8'he6,8'h13,8'hf2,8'h26,8'h9b, \
  8'hbc,8'hb3,8'h54,8'h62,8'h6e,8'h36,8'h13,8'h67, \
  8'h8c,8'hdf,8'hcf,8'hf4,8'hd4,8'h6a,8'h2b,8'h0f, \
  8'hd9,8'h1d,8'h33,8'hbc,8'h74,8'ha9,8'h7d,8'hf2, \
  8'hae,8'h3b,8'h55,8'h19,8'h89,8'h41,8'hff,8'hee, \
  8'h78,8'hc8,8'h90,8'h1c,8'hd9,8'hf3,8'h1d,8'hc2, \
  8'hb0,8'h0e,8'h72,8'h2f,8'h02,8'heb,8'haa,8'h27, \
  8'hbc,8'he9,8'h1b,8'hd8,8'h4a,8'h59,8'hcb,8'hf1, \
  8'h4e,8'h90,8'h00,8'he1,8'hb0,8'h4a,8'h68,8'h78, \
  8'h9d,8'h7c,8'h98,8'h29,8'ha5,8'h6a,8'h7d,8'hee, \
  8'h91,8'h49,8'h3d,8'h61,8'h37,8'hb7,8'h4d,8'h3a, \
  8'he9,8'hdc,8'ha2,8'h52,8'ha9,8'hb9,8'h05,8'h4f, \
  8'h4b,8'h1b,8'h8f,8'h6a,8'h4f,8'hc1,8'h17,8'h57, \
  8'he3,8'ha6,8'hd0,8'h7f,8'h9a,8'h4d,8'hd0,8'h07, \
  8'h5c,8'h44,8'h97,8'h24,8'hfc,8'hf0,8'h95,8'h83, \
  8'h65,8'h51,8'h81,8'h5b,8'h75,8'hde,8'h76,8'h17, \
  8'hfb,8'hea,8'hba,8'h79,8'h5b,8'h1b,8'h6f,8'h21, \
  8'h42,8'he1,8'he1,8'h85,8'h16,8'h69,8'hc0,8'h95, \
  8'haf,8'h48,8'h93,8'h5f,8'he6,8'hc8,8'h32,8'h61, \
  8'hc1,8'hc7,8'h76,8'h73,8'h5d,8'hf2,8'hfb,8'h0a, \
  8'h64,8'hc9,8'h61,8'h7c,8'hb1,8'hbc,8'h4e,8'hdb, \
  8'h88,8'h79,8'h47,8'he6,8'h09,8'hdf,8'h2d,8'h7f, \
  8'h9e,8'h7e,8'hea,8'h88,8'h47,8'hbc,8'h97,8'hbb, \
  8'h5f,8'h7b,8'hc5,8'h45,8'h36,8'hec,8'h25,8'h99, \
  8'h66,8'hf0,8'he0,8'h82,8'ha0,8'ha8,8'h8e,8'ha7, \
  8'h27,8'h3d,8'h50,8'hda,8'hd5,8'h01,8'hdf,8'hb4, \
  8'ha7,8'h4b,8'h28,8'h64,8'hf6,8'h22,8'h59,8'h5c, \
  8'hbf,8'hf3,8'h10,8'h93,8'hc6,8'hcf,8'hda,8'h48, \
  8'hcb,8'hbc,8'hdc,8'h34,8'h80,8'h15,8'h4d,8'h4e, \
  8'hee,8'h4d,8'h36,8'hf8,8'h33,8'he9,8'hf9,8'h46, \
  8'ha1,8'h81,8'h69,8'hcb,8'h72,8'h82,8'hac,8'hd8, \
  8'hdd,8'hf3,8'hec,8'h42,8'hfb,8'hf5,8'h76,8'h8c, \
  8'he7,8'h29,8'h05,8'h00,8'hbb,8'hea,8'h12,8'h56, \
  8'hae,8'h29,8'h0e,8'haf,8'h94,8'haa,8'h99,8'he8, \
  8'h92,8'h22,8'h53,8'hd2,8'h10,8'hf4,8'h2d,8'ha0, \
  8'ha1,8'hac,8'hff,8'h38,8'hb0,8'h00,8'h80,8'h5c, \
  8'h6b,8'h49,8'h93,8'h60,8'haf,8'hc5,8'hb1,8'hb2, \
  8'h63,8'h40,8'h7b,8'hf5,8'hb0,8'hd8,8'ha7,8'hd0, \
  8'hdd,8'ha8,8'h3a,8'h50,8'h16,8'h9b,8'h9c,8'h68, \
  8'h9b,8'he7,8'hd4,8'hf9,8'h79,8'had,8'h84,8'h7b, \
  8'h8f,8'hf5,8'hfe,8'h77,8'hb7,8'he6,8'h08,8'ha1, \
  8'h26,8'haf,8'had,8'h12,8'h62,8'h7c,8'ha9,8'h93, \
  8'h9c,8'h31,8'ha3,8'hb4,8'h22,8'hce,8'h1a,8'h6f, \
  8'h87,8'hf0,8'h05,8'hef,8'h90,8'h01,8'h05,8'h1b, \
  8'h50,8'hde,8'h69,8'h59,8'h62,8'hf9,8'h49,8'hda, \
  8'h79,8'hd8,8'h0b,8'hbf,8'h92,8'h90,8'h55,8'hab, \
  8'he7,8'h50,8'h42,8'h0f,8'h5f,8'hb5,8'h33,8'hd6, \
  8'h96,8'h24,8'ha7,8'hb9,8'hd5,8'h0a,8'hf2,8'h61, \
  8'h25,8'h7f,8'h3e,8'h36,8'h3c,8'ha8,8'h19,8'h78, \
  8'h30,8'h19,8'h14,8'h88,8'hfc,8'h60,8'h91,8'he2, \
  8'h09,8'hea,8'hae,8'hc6,8'h27,8'hf6,8'ha9,8'h83, \
  8'h11,8'h20,8'hbd,8'hea,8'ha7,8'hfe,8'haf,8'h2f, \
  8'hc1,8'hc6,8'h96,8'h17,8'h2b,8'h94,8'ha9,8'h2c, \
  8'h44,8'h6a,8'h2f,8'hcd,8'he3,8'h12,8'h60,8'hc9, \
  8'h99,8'hdb,8'h12,8'hce,8'h97,8'h14,8'h95,8'hd7, \
  8'he6,8'hdb,8'h43,8'h5d,8'h84,8'h50,8'hbf,8'hda, \
  8'h8e,8'hf0,8'he0,8'hfd,8'h18,8'h25,8'h48,8'h32, \
  8'h51,8'hdd,8'he2,8'haa,8'he7,8'hbe,8'hff,8'h3f, \
  8'h53,8'hd4,8'h57,8'hf8,8'h3a,8'hce,8'h83,8'h52, \
  8'h04,8'h11,8'h0c,8'hf2,8'h2b,8'h85,8'h97,8'h39, \
  8'h0b,8'h18,8'hc4,8'h59,8'hb3,8'h31,8'h7d,8'h8c, \
  8'h43,8'hb6,8'h2e,8'h08,8'h9d,8'h7e,8'hae,8'h79, \
  8'h31,8'h24,8'hd6,8'h03,8'h5b,8'h7c,8'h78,8'he9, \
  8'h61,8'he2,8'h3e,8'h2d,8'h29,8'h4d,8'hc4,8'h72, \
  8'hf1,8'h3c,8'h75,8'h17,8'h93,8'hb2,8'hd2,8'h49, \
  8'h1b,8'h9d,8'h43,8'hf7,8'h0c,8'h75,8'hec,8'h03, \
  8'hba,8'h29,8'hcb,8'ha6,8'h65,8'h90,8'hf6,8'h2b, \
  8'h31,8'hb8,8'h98,8'h4c,8'h5b,8'h51,8'h1c,8'h34, \
  8'hc6,8'hf6,8'h2d,8'h7a,8'h8f,8'h92,8'hf1,8'h9f, \
  8'h71,8'h97,8'h07,8'h09,8'hc0,8'hce,8'hb1,8'h6e, \
  8'h53,8'hd3,8'h4c,8'hfa,8'h6c,8'hb7,8'h18,8'h16, \
  8'h9f,8'hf7,8'h5f,8'hf6,8'h69,8'h8a,8'h54,8'hc6, \
  8'hac,8'h02,8'h3b,8'ha1,8'h3c,8'ha5,8'h77,8'h64, \
  8'h2b,8'he5,8'hda,8'hfc,8'h46,8'haa,8'h29,8'h95, \
  8'h00,8'hb3,8'h00,8'heb,8'h94,8'hc9,8'h47,8'h4a, \
  8'hac,8'h79,8'h5d,8'h3c,8'h8b,8'h52,8'h02,8'hf5, \
  8'h4a,8'h8c,8'h53,8'h26,8'hee,8'h1d,8'h51,8'h7a, \
  8'hfb,8'ha8,8'he3,8'h3b,8'hcb,8'h88,8'h36,8'he2, \
  8'ha3,8'h3f,8'ha9,8'hc1,8'h99,8'hf8,8'ha3,8'he9, \
  8'h41,8'he0,8'h7f,8'hd3,8'h31,8'hbd,8'h48,8'h1b, \
  8'h9f,8'h9f,8'h4e,8'h7f,8'h89,8'h8a,8'h3d,8'h6c, \
  8'h96,8'h72,8'h25,8'h6b,8'ha8,8'h43,8'h04,8'hba, \
  8'had,8'h1f,8'hd3,8'h59,8'hb2,8'h1e,8'h7d,8'h56, \
  8'hb5,8'h10,8'h1d,8'hf6,8'h87,8'h0c,8'h8b,8'h86, \
  8'h5f,8'h09,8'h3a,8'h5c,8'h1b,8'h52,8'hfc,8'h83, \
  8'h97,8'h90,8'h9a,8'h25,8'h4d,8'hf1,8'hc4,8'h46, \
  8'hcc,8'h15,8'hca,8'hb0,8'h1d,8'hec,8'hae,8'h55, \
  8'h98,8'h3e,8'ha8,8'ha0,8'h11,8'h53,8'h34,8'hfb, \
  8'hdb,8'hc4,8'h0e,8'h10,8'h5d,8'ha5,8'h34,8'h8a, \
  8'h42,8'h6a,8'h86,8'hb4,8'h6d,8'h54,8'h3d,8'h31, \
  8'hee,8'h99,8'he2,8'he7,8'h41,8'hef,8'h60,8'hb1, \
  8'h20,8'h2c,8'h39,8'h49,8'h91,8'h92,8'h62,8'h36, \
  8'hb7,8'hb6,8'h4c,8'h95,8'haa,8'hc7,8'h44,8'h04, \
  8'h45,8'h17,8'h93,8'h76,8'h7b,8'h3a,8'hb1,8'h68, \
  8'h75,8'h40,8'h64,8'h9d,8'h46,8'h39,8'h7d,8'h19, \
  8'h7b,8'hc7,8'h05,8'ha6,8'h1e,8'hc6,8'h50,8'h39, \
  8'h9e,8'h4c,8'h2c,8'h25,8'h1f,8'h7c,8'h2e,8'hfc, \
  8'h5f,8'h7c,8'ha0,8'h8d,8'h53,8'h82,8'hd3,8'h1c, \
  8'h04,8'hef,8'h88,8'hfb,8'h47,8'hd9,8'h56,8'had, \
  8'h0d,8'hdb,8'h45,8'h07,8'ha7,8'ha6,8'h3b,8'h44, \
  8'h52,8'ha4,8'h26,8'h3a,8'hcb,8'h76,8'h47,8'h10, \
  8'h60,8'h39,8'had,8'h9b,8'h6d,8'h12,8'hdd,8'h99, \
  8'h8d,8'h24,8'h45,8'h5a,8'h04,8'h97,8'h1d,8'h36, \
  8'hd1,8'h65,8'haa,8'h7d,8'h17,8'hbd,8'h77,8'h85, \
  8'h0d,8'h68,8'h79,8'hfb,8'ha8,8'hd1,8'h4c,8'hb9, \
  8'hb4,8'h2f,8'hc4,8'hdb,8'h3c,8'h7e,8'h07,8'he7, \
  8'hc0,8'h8e,8'h5b,8'hee,8'h5d,8'h7d,8'h28,8'hfd, \
  8'h23,8'hee,8'h2a,8'h4c,8'h35,8'h55,8'h79,8'hd8, \
  8'h0b,8'h99,8'h91,8'ha7,8'hf4,8'hd3,8'h00,8'h0e, \
  8'h65,8'h44,8'h52,8'hf8,8'h3d,8'h54,8'h3c,8'h17, \
  8'h5a,8'h68,8'ha5,8'h50,8'h23,8'h8f,8'hf9,8'h9c, \
  8'ha4,8'hc2,8'hf8,8'h8a,8'h99,8'h3a,8'h5c,8'hfa, \
  8'hb6,8'h13,8'h89,8'hb1,8'h38,8'h0f,8'h2b,8'hd9, \
  8'h5f,8'hfb,8'ha4,8'h6c,8'h75,8'h19,8'he1,8'he7, \
  8'h7b,8'h92,8'hd9,8'hce,8'h93,8'h63,8'h0d,8'h5a, \
  8'h75,8'h5e,8'ha8,8'hf2,8'h2e,8'h6c,8'h82,8'hb6, \
  8'h52,8'hb4,8'h3f,8'h5c,8'hb9,8'hf8,8'h41,8'hc1, \
  8'hc2,8'hac,8'hca,8'h1f,8'h52,8'hbb,8'h26,8'h76, \
  8'h27,8'h6b,8'h3f,8'ha2,8'h89,8'hd3,8'h63,8'h02, \
  8'hc5,8'h15,8'hb6,8'hcc,8'h7b,8'h08,8'h23,8'h51, \
  8'h43,8'h39,8'h77,8'hec,8'h96,8'hfe,8'he0,8'h56, \
  8'hd2,8'h1b,8'h12,8'h57,8'h9f,8'hfc,8'hb3,8'h2c, \
  8'hb4,8'h86,8'h4d,8'hb6,8'h93,8'h87,8'hec,8'he6, \
  8'h15,8'h71,8'hcc,8'h53,8'haf,8'h0b,8'h20,8'h1d, \
  8'hce,8'h06,8'hb2,8'h48,8'h67,8'hb8,8'hea,8'h38, \
  8'hd2,8'hb9,8'he2,8'hb1,8'h9a,8'h63,8'h6d,8'h3f, \
  8'haa,8'h01,8'hff,8'h9d,8'h6b,8'h4d,8'h92,8'hb6, \
  8'h29,8'hcb,8'h87,8'hf0,8'h71,8'h5b,8'h1c,8'h00, \
  8'hc9,8'h52,8'h66,8'h94,8'h17,8'hcd,8'h95,8'h15, \
  8'h71,8'h88,8'h40,8'hc1,8'h57,8'h5e,8'h77,8'h2f, \
  8'hc1,8'h91,8'h65,8'h6a,8'hb0,8'h7c,8'h61,8'h3f, \
  8'h93,8'he6,8'hf7,8'hab,8'h8e,8'h2b,8'hd8,8'h10, \
  8'hef,8'h1f,8'h1d,8'h81,8'hb9,8'hf1,8'hc1,8'h11, \
  8'hd6,8'hdb,8'h38,8'h62,8'h0d,8'h56,8'h0a,8'h7e, \
  8'hb6,8'h51,8'h91,8'hb2,8'h70,8'he0,8'h56,8'h2f, \
  8'h96,8'h53,8'h6c,8'h33,8'h87,8'h4a,8'ha8,8'h25, \
  8'hab,8'h44,8'hd9,8'h99,8'h6c,8'h89,8'h9a,8'ha5, \
  8'hd9,8'h3e,8'h90,8'h2e,8'h7f,8'h88,8'h5c,8'h94, \
  8'h8c,8'h90,8'hf2,8'h2a,8'hd7,8'hcd,8'hc8,8'h34, \
  8'hf8,8'h24,8'h47,8'h5e,8'h93,8'h21,8'h73,8'h45, \
  8'h6b,8'h65,8'h4d,8'h00,8'h11,8'h54,8'he7,8'hbc, \
  8'h2e,8'h30,8'h9d,8'he7,8'h39,8'h42,8'h64,8'hd1, \
  8'he8,8'h0e,8'h80,8'hd6,8'h92,8'hb2,8'h25,8'hcf, \
  8'h0a,8'h5f,8'he2,8'h94,8'h19,8'h98,8'h12,8'h23, \
  8'hcc,8'h3a,8'hbb,8'h6a,8'he3,8'h66,8'hd4,8'h41, \
  8'h2c,8'hd6,8'h10,8'hde,8'h16,8'hc8,8'h51,8'h6e, \
  8'hda,8'h95,8'h11,8'hd8,8'hf1,8'h53,8'h78,8'ha4, \
  8'hb9,8'h2d,8'h8d,8'hcc,8'h20,8'h17,8'hef,8'h19, \
  8'h0e,8'h4d,8'hcf,8'h45,8'hde,8'hc3,8'hc4,8'h81, \
  8'h01,8'h6b,8'hae,8'h02,8'hd9,8'ha3,8'h2f,8'h95, \
  8'h78,8'h09,8'ha4,8'h11,8'h77,8'h0f,8'h29,8'h49, \
  8'h8a,8'h96,8'h79,8'hf7,8'h4b,8'ha5,8'hae,8'h3b, \
  8'h05,8'hdc,8'hd6,8'h7e,8'hfe,8'ha4,8'h5c,8'hdf, \
  8'h36,8'h66,8'h75,8'hb1,8'ha0,8'h19,8'hd4,8'he4, \
  8'h4d,8'h82,8'h07,8'ha1,8'h01,8'h1f,8'h06,8'h08, \
  8'hb1,8'h31,8'h7f,8'hdc,8'he7,8'h99,8'h88,8'h8d, \
  8'h52,8'he8,8'h26,8'h50,8'hab,8'h85,8'h5d,8'h13, \
  8'h9a,8'h0f,8'h11,8'h9b,8'h99,8'h59,8'hab,8'h4c, \
  8'h5c,8'hdc,8'he4,8'hd1,8'h21,8'hd9,8'h69,8'hc5, \
  8'h02,8'he9,8'h2d,8'h28,8'hc1,8'hf5,8'h76,8'he4, \
  8'h20,8'h4c,8'h7e,8'h9b,8'h9f,8'h5e,8'h5b,8'hd8, \
  8'h9d,8'h3d,8'h3c,8'h08,8'h74,8'h9d,8'h7f,8'h1c, \
  8'he7,8'h8a,8'h88,8'h7a,8'h5a,8'he0,8'h82,8'hff, \
  8'h11,8'hea,8'hc5,8'hbd,8'h7a,8'ha8,8'h1e,8'haa, \
  8'h19,8'h79,8'h4c,8'h25,8'hb1,8'h91,8'hd0,8'hab, \
  8'hd6,8'h31,8'h4f,8'h1d,8'h59,8'h1e,8'h21,8'hec, \
  8'hcf,8'h58,8'hfb,8'h5b,8'hab,8'h4f,8'heb,8'h44, \
  8'hf0,8'h96,8'h4e,8'h6c,8'hf7,8'h45,8'h48,8'h22, \
  8'ha9,8'h5b,8'hea,8'h50,8'hfa,8'h8c,8'h79,8'hf5, \
  8'h64,8'h8a,8'h30,8'hc6,8'h63,8'hf9,8'hf9,8'h72, \
  8'h5d,8'h91,8'h2a,8'hef,8'h81,8'h5a,8'hde,8'hcc, \
  8'h08,8'h5b,8'h15,8'h06,8'hd3,8'h4e,8'h18,8'h0d, \
  8'h89,8'h94,8'h25,8'h0c,8'h03,8'h64,8'h34,8'ha4, \
  8'hd6,8'hd3,8'hb7,8'ha6,8'h41,8'h98,8'h42,8'hb5, \
  8'h7e,8'hd4,8'h66,8'h64,8'ha7,8'h92,8'hb1,8'h55, \
  8'h1c,8'hba,8'h81,8'h7e,8'ha9,8'hf3,8'hda,8'ha9, \
  8'h69,8'hcc,8'h28,8'h55,8'h67,8'hd8,8'hed,8'h98, \
  8'h82,8'h99,8'h61,8'had,8'h67,8'h9a,8'h03,8'hbd, \
  8'h92,8'hde,8'hd9,8'hfb,8'h23,8'hf0,8'h69,8'hd3, \
  8'hda,8'hac,8'hc5,8'h28,8'h02,8'hb5,8'h3e,8'h29, \
  8'h23,8'h47,8'h13,8'h7d,8'hcf,8'h3d,8'h9a,8'h48, \
  8'hc1,8'h23,8'h5e,8'h68,8'hb0,8'h9c,8'h0b,8'hbc, \
  8'h4d,8'hc8,8'hab,8'h3f,8'had,8'hed,8'hdd,8'hc5, \
  8'h89,8'hc1,8'h00,8'hf3,8'hc8,8'he7,8'hd5,8'h11, \
  8'h5a,8'h28,8'hf7,8'h88,8'h21,8'h94,8'hbf,8'h85, \
  8'h56,8'hf7,8'hfa,8'h7b,8'h19,8'h57,8'hcb,8'h87, \
  8'h93,8'hfb,8'h0b,8'heb,8'h8e,8'h1b,8'h3c,8'h5b, \
  8'ha4,8'h08,8'h61,8'haa,8'ha8,8'h7a,8'h1e,8'hdf, \
  8'heb,8'h62,8'hc6,8'hde,8'hfe,8'hb7,8'h65,8'hb6, \
  8'ha3,8'h90,8'he8,8'h3e,8'h9b,8'h0e,8'hba,8'h61, \
  8'ha3,8'h56,8'h25,8'hfc,8'hb2,8'h99,8'h27,8'h70, \
  8'he7,8'h3f,8'hce,8'heb,8'h82,8'h55,8'hb2,8'hdf, \
  8'h4f,8'he9,8'hdb,8'h57,8'h20,8'hc2,8'h34,8'h64, \
  8'h33,8'h26,8'hc3,8'hfc,8'h7d,8'ha5,8'ha6,8'h77, \
  8'h68,8'ha3,8'h55,8'hbf,8'hb9,8'hf0,8'h7b,8'h85, \
  8'ha9,8'hf4,8'hcf,8'h0d,8'h93,8'h08,8'hc6,8'he7, \
  8'hd3,8'hdd,8'h29,8'hca,8'h7a,8'h11,8'h0c,8'hbf, \
  8'h81,8'h65,8'h96,8'h7f,8'h88,8'ha3,8'h5e,8'h95, \
  8'h15,8'h5a,8'h26,8'h2d,8'had,8'h7b,8'hc4,8'h6c, \
  8'hfd,8'h88,8'hed,8'h23,8'hdd,8'hb0,8'h0b,8'hcc, \
  8'hb5,8'h09,8'h02,8'hd2,8'h96,8'h1e,8'h36,8'h68, \
  8'h52,8'h4d,8'h7f,8'hc6,8'hf2,8'h64,8'h73,8'h24, \
  8'h7f,8'h88,8'hea,8'h56,8'h23,8'h1b,8'h75,8'h64, \
  8'h4a,8'ha7,8'hfe,8'h7b,8'h97,8'h63,8'he9,8'h88, \
  8'h7b,8'h7d,8'h91,8'h7a,8'hde,8'hf1,8'h52,8'h85, \
  8'h27,8'hf6,8'h5a,8'h57,8'h7d,8'h7e,8'hae,8'h0b, \
  8'h06,8'h08,8'h56,8'h67,8'h2f,8'h54,8'h2b,8'hda, \
  8'h24,8'hec,8'had,8'h4f,8'h34,8'h11,8'h05,8'hbf, \
  8'h67,8'hb1,8'hdc,8'h0e,8'h8a,8'h64,8'ha1,8'hea, \
  8'hbe,8'h67,8'h5a,8'he5,8'h5c,8'haa,8'h97,8'h18, \
  8'h5f,8'h9a,8'h24,8'h86,8'h7f,8'h17,8'hb9,8'hac, \
  8'h4e,8'h77,8'h48,8'hba,8'h32,8'h32,8'h07,8'h36, \
  8'hda,8'h95,8'h2c,8'hdb,8'hde,8'hfb,8'h11,8'h13, \
  8'ha8,8'hd4,8'he4,8'h1e,8'hcb,8'h8b,8'hc9,8'h68, \
  8'hb6,8'he0,8'hb5,8'h7d,8'h15,8'hf7,8'h75,8'h71, \
  8'h98,8'h37,8'h2e,8'h85,8'h28,8'h32,8'hc3,8'h83, \
  8'h7b,8'h2a,8'h3a,8'h34,8'h2d,8'h04,8'h18,8'h31, \
  8'hab,8'h0f,8'hdb,8'h7b,8'h7f,8'h2a,8'h29,8'hcb, \
  8'h32,8'h52,8'h2e,8'h55,8'h88,8'hc0,8'h0a,8'h41, \
  8'he6,8'h2d,8'h7b,8'h48,8'hf2,8'hc8,8'h52,8'h16, \
  8'h0f,8'hed,8'h80,8'he6,8'hb8,8'hb3,8'hac,8'h94 \
  }
